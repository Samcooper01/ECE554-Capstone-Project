module MEMORY_STORE(iFRAMECOUNT, iDVAL, iGray, oGray, oDVAL);
    // Inputs
    input [31:0] iFRAMECOUNT;
    input iDVAL;
    input [11:0] iGray;
    
    // Outputs
    output oGray;
    output oDVAL;







endmodule