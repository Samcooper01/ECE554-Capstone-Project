// Top level file for everything